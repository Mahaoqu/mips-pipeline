`timescale 1ns / 1ps
module SoC(input clk, input rst);
    SoC_design soc(.clk(clk), .rst(rst));
endmodule